module MOD14_counter(
    input clk,
    output ff0,
    output ff1,
    output ff2,
    output ff3
);

    

endmodule