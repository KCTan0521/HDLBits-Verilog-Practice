module top_module(
	input clk, 
	input load, 
	input [9:0] data, 
	output tc
);

    reg [9:0] counter;

    always @(posedge clk) begin
        if (load) begin
            counter <= data;
        end
        else begin
            if (counter > 0 ) begin
                counter <= counter - 1'b1;
            end
            else begin
                counter <= 1'b0;
            end
        end
    end

    assign tc = counter == 10'b0;
endmodule
